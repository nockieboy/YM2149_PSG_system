/************************************************************************************************************************************* 

This DAC LUT table was created with the 'BHG_jt49_exp_tablegen.v', v1.0, Aug 6, 2022.
                                         It was rendered using Modelsim.
                                         by Brian Guralnick.
                                         https://github.com/BrianHGinc

Table generated using a LSB_DB_CORRECTION setting of [8:12] :'{ 15, 14, 13, 12, 11}.
                                                              *** 15 is optimum for an 8 bit dac ***.

This code is free to use.  Just be fair and give credit where it is due.

******************************************************************
*** This code was written by BrianHG providing an optional     ***
*** volume decibel attenuation with taper optimization for     ***
*** the first few DAC volume steps.                            ***
*** This code will generate LUT tables for 8 to 12 bit DACs.   ***
******************************************************************/

// *************************************************************************************************************************************
// *** 8  bit DAC LUT with a dynamic range of -48 decibels.
// *************************************************************************************************************************************
localparam logic [15:0] dlut_8  [0:31] = '{   0,   1,   2,   3,   4,   5,   6,   8,  10,  12,  14,  17,  19,  23,  26,  31,
                                             35,  41,  47,  54,  62,  70,  80,  92, 104, 119, 135, 154, 175, 198, 225, 255};
// *************************************************************************************************************************************
// *** 9  bit DAC LUT with a dynamic range of -54 decibels.
// *************************************************************************************************************************************
localparam logic [15:0] dlut_9  [0:31] = '{   0,   1,   2,   3,   4,   6,   7,   9,  12,  14,  17,  21,  25,  30,  36,  42,
                                             50,  59,  69,  81,  95, 111, 130, 151, 177, 206, 240, 279, 325, 378, 439, 511};
// *************************************************************************************************************************************
// *** 10 bit DAC LUT with a dynamic range of -60 decibels.
// *************************************************************************************************************************************
localparam logic [15:0] dlut_10 [0:31] = '{   0,   1,   2,   3,   5,   6,   8,  11,  14,  17,  21,  26,  32,  39,  48,  58,
                                             70,  84, 101, 121, 145, 174, 208, 248, 297, 354, 423, 505, 603, 719, 858,1023};
// *************************************************************************************************************************************
// *** 11 bit DAC LUT with a dynamic range of -66 decibels.
// *************************************************************************************************************************************
localparam logic [15:0] dlut_11 [0:31] = '{   0,   1,   2,   3,   5,   7,   9,  12,  16,  20,  26,  33,  41,  51,  63,  78,
                                             96, 118, 146, 179, 220, 270, 331, 406, 497, 609, 745, 913,1117,1367,1673,2047};
// *************************************************************************************************************************************
// *** 12 bit DAC LUT with a dynamic range of -72 decibels.
// *************************************************************************************************************************************
localparam logic [15:0] dlut_12 [0:31] = '{   0,   1,   2,   3,   5,   8,  10,  14,  18,  24,  31,  40,  51,  65,  82, 104,
                                            132, 166, 209, 264, 332, 418, 526, 661, 830,1043,1311,1647,2068,2597,3261,4095};

// **********************************************
// *** Coalesce the 5 tables into a 2D array. ***
// **********************************************
localparam logic [15:0] dlut_sel [8:12][0:31] = '{ dlut_8, dlut_9, dlut_10, dlut_11, dlut_12 };

// *** Table End.

